`ifndef LWC_CONSTANTS_VH
`define LWC_CONSTANTS_VH

parameter ASYNC_RSTN = 1;

`endif