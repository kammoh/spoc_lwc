parameter ASYNC_RSTN = 1;